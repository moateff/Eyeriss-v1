package cfg_pkg;
import shared_pkg::*;
    
    task conv1_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/conv1/serial_data.txt";
        cfg_scan_chain(filename);
    endtask
    
    task conv2_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/conv2/serial_data.txt";
        cfg_scan_chain(filename);
    endtask
    
    task conv3_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/conv3/serial_data.txt";
        cfg_scan_chain(filename);
    endtask
    
    task conv4_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/conv4/serial_data.txt";
        cfg_scan_chain(filename);
    endtask
    
    task conv5_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/conv5/serial_data.txt";
        cfg_scan_chain(filename);
    endtask

    task max1_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/max1/serial_data.txt";
        cfg_scan_chain(filename);
    endtask

    task max2_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/max2/serial_data.txt";
        cfg_scan_chain(filename);
    endtask
            
    task max3_cfg();
        string filename;
        filename = "D:/data/Graduation Project/GP_AlexNet/WE Scan Chain/sw/max3/serial_data.txt";
        cfg_scan_chain(filename);
    endtask  
      
    task cfg_scan_chain(
        input string filename
    );
        int file;
        int char_val;
        int bit_val;
        string line;

        file = $fopen(filename, "r");
        if (file == 0) begin
            $display("[ERROR] Could not open file: %s", filename);
            $stop;
        end

        shared_pkg::scan_enable = 1;

        while (!$feof(file)) begin
            line = "";
            void'($fgets(line, file));
            if (line.len() > 0) begin
            $sscanf(line, "%d", bit_val);
            shared_pkg::scan_in = bit_val;
            wait_link_cycle(1);
            end
        end

        shared_pkg::scan_enable = 0;
        $fclose(file);

    endtask
    
    /*
    int expected_q_enable       [0:11][0:13]; 
    int expected_q_LN_sel       [0:11][0:13]; 
    int expected_ifmap_row_ids  [0:11];
    int expected_ifmap_col_ids  [0:11][0:13];
    int expected_filter_row_ids [0:11];
    int expected_filter_col_ids [0:11][0:13];
    int expected_ipsum_row_ids  [0:11];
    int expected_ipsum_col_ids  [0:11][0:13];
    int expected_opsum_row_ids  [0:11];
    int expected_opsum_col_ids  [0:11][0:13];
    
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/serial_data.txt"; //directory of the file generated by the script
    configure_scan_chain(filename);
    
    wait_core_cycle(3500);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/parameters.txt";
    check_parameters_from_file (filename);

    wait_core_cycle(1);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/enables.txt";
    read_q_enable_file(filename);

    wait_core_cycle(1);
    check_q_enable_with_dut();

    wait_core_cycle(1);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/ln_selectors.txt";
    read_q_LN_sel_file(filename);

    wait_core_cycle(1);
    check_q_LN_sel_with_dut();*
    wait_core_cycle(3500);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/ifmap_ids.txt";
    read_matrix_file(filename,expected_ifmap_row_ids,expected_ifmap_col_ids);
    
    wait_core_cycle(1);
    compare_ifmap_ids(expected_ifmap_row_ids,expected_ifmap_col_ids);
    
    
    wait_core_cycle(3500);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/filters_ids.txt";
    read_matrix_file(filename,expected_filter_row_ids,expected_filter_col_ids);
    
    wait_core_cycle(1);
    compare_ifmap_ids(expected_filter_row_ids,expected_filter_col_ids);*
    wait_core_cycle(3500);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/ipsum_ids.txt";
    read_matrix_file(filename,expected_ipsum_row_ids,expected_ipsum_col_ids);
    
    wait_core_cycle(1);
    compare_ifmap_ids(expected_ipsum_row_ids,expected_ipsum_col_ids);
    *
    wait_core_cycle(1);
    filename = "E:/9th10th GP/GP_AlexNet/WE Scan Chain/sw/conv1/opsum_ids.txt";
    read_matrix_file(filename,expected_opsum_row_ids,expected_opsum_col_ids);
    
    wait_core_cycle(1);
    compare_ifmap_ids(expected_opsum_row_ids,expected_opsum_col_ids);

    task read_q_enable_file(input string filename);
        int file, r, c;
        int val;
        begin
            file = $fopen(filename, "r");
            if (file == 0) begin
                $display("ERROR: Cannot open file: %s", filename);
                $finish;
            end

            r = 0;
            while (!$feof(file) && r < 12) begin
                for (c = 0; c < 14; c++) begin
                    $fscanf(file, "%d", val);
                    expected_q_enable[r][c] = val;
                end
                r++;
            end

            $fclose(file);
            $display("Enables loaded into expected_q_enable[][]");
        end
    endtask

    task read_q_LN_sel_file(input string filename);
        int file, r, c;
        int val, status;
        begin
            file = $fopen(filename, "r");
            if (file == 0) begin
                $display("ERROR: Cannot open file: %s", filename);
                $finish;
            end

            r = 0;
            while (!$feof(file) && r < 12) begin
                for (c = 0; c < 14; c++) begin
                    status = $fscanf(file, "%d", val);
                    if (status != 1) begin
                        $display("WARNING: Invalid data at r=%0d, c=%0d", r, c);
                        val = 0; // or some default
                    end
                    expected_q_LN_sel[r][c] = val;
                end
                r++;
            end

            $fclose(file);
            $display("ln_selectors.txt loaded into expected_q_LN_sel[][]");
        end
    endtask

    task read_matrix_file(
        input  string filename,
        output int    row_ids [0:11],        // 12 rows
        output int    col_ids [0:11][0:13]   // 12 rows � 14 cols
    );
        int file, status;
        int r, c, temp;

        begin
            file = $fopen(filename, "r");
            if (file == 0) begin
                $display("[ERROR] Cannot open file: %s", filename);
                $finish;
            end

            for (r = 0; r < 12; r++) begin
                // Read row ID (first column)
                status = $fscanf(file, "%d", temp);
                if (status != 1) begin
                    $display("[ERROR] Failed to read row ID at row %0d", r);
                    $finish;
                end
                row_ids[r] = temp;

                // Read col IDs (remaining 14 columns)
                for (c = 0; c < 14; c++) begin
                    status = $fscanf(file, "%d", temp);
                    if (status != 1) begin
                        $display("[ERROR] Failed to read col ID at row %0d, col %0d", r, c);
                        $finish;
                    end
                    col_ids[r][c] = temp;
                end
            end

            $fclose(file);
            $display("[INFO] Successfully read matrix file: %s", filename);
        end
    endtask

    task compare_signal(input string param_name, input int actual, input int expected);
        if (actual !== expected)
            $display("%s [Mismatch] expected %0d, got %0d", param_name, expected, actual);
    endtask
    
    task check_parameters_from_file(input string filename);
        int file, expected_val;
        string line, name;

        begin
            file = $fopen(filename, "r");
            if (file == 0) begin
            $display("ERROR: Could not open parameter file: %s", filename);
            $finish;
            end

            $display("=== Checking Parameters from %s ===", filename);
            while (!$feof(file)) begin
            line = "";
            void'($fgets(line, file));
            if (line.len() > 0) begin
                $sscanf(line, "%s = %d", name, expected_val);

                // Compare each known parameter name
                if (name == "H")  compare_signal("H", DUT.PARAMETERS.H, expected_val);
                else if (name == "R")  compare_signal("R", DUT.PARAMETERS.R, expected_val);
                else if (name == "E")  compare_signal("E", DUT.PARAMETERS.E, expected_val);
                else if (name == "C")  compare_signal("C", DUT.PARAMETERS.C, expected_val);
                else if (name == "M")  compare_signal("M", DUT.PARAMETERS.M, expected_val);
                else if (name == "N")  compare_signal("N", DUT.PARAMETERS.N, expected_val);
                else if (name == "U")  compare_signal("U", DUT.PARAMETERS.U, expected_val);
                else if (name == "V")  compare_signal("V", DUT.PARAMETERS.V, expected_val);
                else if (name == "n")  compare_signal("n", DUT.PARAMETERS.n, expected_val);
                else if (name == "e")  compare_signal("e", DUT.PARAMETERS.e, expected_val);
                else if (name == "p")  compare_signal("p", DUT.PARAMETERS.p, expected_val);
                else if (name == "q")  compare_signal("q", DUT.PARAMETERS.q, expected_val);
                else if (name == "r")  compare_signal("r", DUT.PARAMETERS.r, expected_val);
                else if (name == "t")  compare_signal("t", DUT.PARAMETERS.t, expected_val);
                else if (name == "X")  compare_signal("X", DUT.PARAMETERS.X, expected_val);
                else
                $display("Unknown parameter: %s", name);
            end
            end
            $fclose(file);
             $display("=== Checking Parameters Finished  ===");
        end
    endtask
    
    task check_q_enable_with_dut;
        int r, c;
        bit dut_val, expected_val;
        automatic int mismatch_count = 0;
        
        begin
            $display("=== Comparing q_enable[][] with expected values ===");
            for (r = 0; r < 12; r++) begin
                for (c = 0; c < 14; c++) begin
                    expected_val = expected_q_enable[r][c];
                    dut_val = DUT.PROCESSING.pe_array_inst.pe_array_inst.enable[r][c];

                    if (dut_val !== expected_val) begin
                        $display("[Mismatch] at q_enable[%0d][%0d]: DUT=%0b, Expected=%0b", r, c, dut_val, expected_val);
                        mismatch_count++;
                    end
                end
            end
            $display("=== Comparison Finished: %0d mismatches found ===", mismatch_count);
        end
    endtask

    task check_q_LN_sel_with_dut;
        int r, c;
        bit dut_val, expected_val;
        automatic int mismatch_count = 0;
        begin
            $display("=== Comparing q_LN_sel[][] with expected values ===");
            for (r = 0; r < 12; r++) begin
                for (c = 0; c < 14; c++) begin
                    expected_val = expected_q_LN_sel[r][c];
                    dut_val = DUT.PROCESSING.pe_array_inst.pe_array_inst.ln_sel[r][c];
    
                    if (dut_val !== expected_val) begin
                    $display("[Mismatch] at q_LN_sel[%0d][%0d]: DUT=%0b, Expected=%0b", r, c, dut_val, expected_val);
                    mismatch_count++;
                end
            end
            end
            $display("=== Comparison Finished: %0d mismatches found ===", mismatch_count);
        end
    endtask
    
    function int get_dut_row_id(input int r);
        case (r)
            0 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0 ].mcc_inst.q_id;
            1 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1 ].mcc_inst.q_id;
            2 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2 ].mcc_inst.q_id;
            3 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3 ].mcc_inst.q_id;
            4 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4 ].mcc_inst.q_id;
            5 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5 ].mcc_inst.q_id;
            6 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6 ].mcc_inst.q_id;
            7 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7 ].mcc_inst.q_id;
            8 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8 ].mcc_inst.q_id;
            9 : get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9 ].mcc_inst.q_id;
            10: get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].mcc_inst.q_id;
            11: get_dut_row_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].mcc_inst.q_id;
            default: begin
                get_dut_row_id = -1;
                $display("[ERROR] Invalid row index: %0d", r);
            end
        endcase
    endfunction

    function int get_dut_col_id(input int r, input int c);
            case (r)
                0: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[0].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                1: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[1].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                2: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[2].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                3: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[3].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                4: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[4].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                5: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[5].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                6: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[6].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                7: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[7].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                8: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[8].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                9: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[9].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                10: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[10].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                11: case (c)
                    0 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[0].mcc_inst.q_id;
                    1 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[1].mcc_inst.q_id;
                    2 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[2].mcc_inst.q_id;
                    3 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[3].mcc_inst.q_id;
                    4 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[4].mcc_inst.q_id;
                    5 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[5].mcc_inst.q_id;
                    6 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[6].mcc_inst.q_id;
                    7 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[7].mcc_inst.q_id;
                    8 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[8].mcc_inst.q_id;
                    9 : get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[9].mcc_inst.q_id;
                    10: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[10].mcc_inst.q_id;
                    11: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[11].mcc_inst.q_id;
                    12: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[12].mcc_inst.q_id;
                    13: get_dut_col_id = eyeriss_tb.DUT.PROCESSING.pe_array_inst.pe_array_inst.ipsum_gin_inst.gin_inst.ROW_MCC_XBUS[11].xbus_inst.MCC_INSTANCE[13].mcc_inst.q_id;
                    default: get_dut_col_id = -1;
                endcase
                default: get_dut_col_id = -1;
            endcase
    endfunction
    
    task compare_ifmap_ids(
        input int row_ids   [0:11],
        input int col_ids   [0:11][0:13]
    );
        
        int dut_row_val, dut_col_val;
        int r, c;
        automatic bit mismatch = 0;

        $display("=== Comparing IDs with DUT ===");
        
            for (r = 0; r < 12; r++) begin
                // Compare row ID
                dut_row_val = get_dut_row_id(r);
                //$display("q_id = %0d",dut_row_val);
                if (row_ids[r] !== dut_row_val) begin
                    $display("[Mismatch][Row %0d] ROW_ID: Expected = %0d, DUT = %0d", r, row_ids[r], dut_row_val);
                    mismatch = 1;
                end

                // Compare col IDs
                for (c = 0; c < 14; c++) begin
                    dut_col_val = get_dut_col_id(r, c);
                    //$display("q_id = %0d",dut_col_val);
                    if (col_ids[r][c] !== dut_col_val) begin
                        $display("[Mismatch][Row %0d, Col %0d] COL_ID: Expected = %0d, DUT = %0d", r, c, col_ids[r][c], dut_col_val);
                        mismatch = 1;
                    end
                end
            end

            if (!mismatch)
                $display("[PASS] All OPSUM_IDS values matched with DUT.");
            else
                $display("[FAIL] One or more OPSUM_IDS values mismatched.");
    endtask
    */
endpackage : cfg_pkg